module analog_top (

);
endmodule