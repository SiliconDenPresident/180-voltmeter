module digital_top (

);

endmodule